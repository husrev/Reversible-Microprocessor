`timescale 1ns / 1ps
	module encoder8_12(
	input [7:0] data_in,
	output reg [11:0] data_out
);
always @*
case(data_in)
	8'b00000000:  data_out <= 12'b000000000000;
	8'b00000001:  data_out <= 12'b000000000111;
	8'b00000010:  data_out <= 12'b000000011001;
	8'b00000011:  data_out <= 12'b000000011110;
	8'b00000100:  data_out <= 12'b000000101010;
	8'b00000101:  data_out <= 12'b000000101101;
	8'b00000110:  data_out <= 12'b000000110011;
	8'b00000111:  data_out <= 12'b000000110100;
	8'b00001000:  data_out <= 12'b000001001011;
	8'b00001001:  data_out <= 12'b000001001100;
	8'b00001010:  data_out <= 12'b000001010010;
	8'b00001011:  data_out <= 12'b000001010101;
	8'b00001100:  data_out <= 12'b000001100001;
	8'b00001101:  data_out <= 12'b000001100110;
	8'b00001110:  data_out <= 12'b000001111000;
	8'b00001111:  data_out <= 12'b000001111111;
	8'b00010000:  data_out <= 12'b000110000001;
	8'b00010001:  data_out <= 12'b000110000110;
	8'b00010010:  data_out <= 12'b000110011000;
	8'b00010011:  data_out <= 12'b000110011111;
	8'b00010100:  data_out <= 12'b000110101011;
	8'b00010101:  data_out <= 12'b000110101100;
	8'b00010110:  data_out <= 12'b000110110010;
	8'b00010111:  data_out <= 12'b000110110101;
	8'b00011000:  data_out <= 12'b000111001010;
	8'b00011001:  data_out <= 12'b000111001101;
	8'b00011010:  data_out <= 12'b000111010011;
	8'b00011011:  data_out <= 12'b000111010100;
	8'b00011100:  data_out <= 12'b000111100000;
	8'b00011101:  data_out <= 12'b000111100111;
	8'b00011110:  data_out <= 12'b000111111001;
	8'b00011111:  data_out <= 12'b000111111110;
	8'b00100000:  data_out <= 12'b001010000010;
	8'b00100001:  data_out <= 12'b001010000101;
	8'b00100010:  data_out <= 12'b001010011011;
	8'b00100011:  data_out <= 12'b001010011100;
	8'b00100100:  data_out <= 12'b001010101000;
	8'b00100101:  data_out <= 12'b001010101111;
	8'b00100110:  data_out <= 12'b001010110001;
	8'b00100111:  data_out <= 12'b001010110110;
	8'b00101000:  data_out <= 12'b001011001001;
	8'b00101001:  data_out <= 12'b001011001110;
	8'b00101010:  data_out <= 12'b001011010000;
	8'b00101011:  data_out <= 12'b001011010111;
	8'b00101100:  data_out <= 12'b001011100011;
	8'b00101101:  data_out <= 12'b001011100100;
	8'b00101110:  data_out <= 12'b001011111010;
	8'b00101111:  data_out <= 12'b001011111101;
	8'b00110000:  data_out <= 12'b001100000011;
	8'b00110001:  data_out <= 12'b001100000100;
	8'b00110010:  data_out <= 12'b001100011010;
	8'b00110011:  data_out <= 12'b001100011101;
	8'b00110100:  data_out <= 12'b001100101001;
	8'b00110101:  data_out <= 12'b001100101110;
	8'b00110110:  data_out <= 12'b001100110000;
	8'b00110111:  data_out <= 12'b001100110111;
	8'b00111000:  data_out <= 12'b001101001000;
	8'b00111001:  data_out <= 12'b001101001111;
	8'b00111010:  data_out <= 12'b001101010001;
	8'b00111011:  data_out <= 12'b001101010110;
	8'b00111100:  data_out <= 12'b001101100010;
	8'b00111101:  data_out <= 12'b001101100101;
	8'b00111110:  data_out <= 12'b001101111011;
	8'b00111111:  data_out <= 12'b001101111100;
	8'b01000000:  data_out <= 12'b010010000011;
	8'b01000001:  data_out <= 12'b010010000100;
	8'b01000010:  data_out <= 12'b010010011010;
	8'b01000011:  data_out <= 12'b010010011101;
	8'b01000100:  data_out <= 12'b010010101001;
	8'b01000101:  data_out <= 12'b010010101110;
	8'b01000110:  data_out <= 12'b010010110000;
	8'b01000111:  data_out <= 12'b010010110111;
	8'b01001000:  data_out <= 12'b010011001000;
	8'b01001001:  data_out <= 12'b010011001111;
	8'b01001010:  data_out <= 12'b010011010001;
	8'b01001011:  data_out <= 12'b010011010110;
	8'b01001100:  data_out <= 12'b010011100010;
	8'b01001101:  data_out <= 12'b010011100101;
	8'b01001110:  data_out <= 12'b010011111011;
	8'b01001111:  data_out <= 12'b010011111100;
	8'b01010000:  data_out <= 12'b010100000010;
	8'b01010001:  data_out <= 12'b010100000101;
	8'b01010010:  data_out <= 12'b010100011011;
	8'b01010011:  data_out <= 12'b010100011100;
	8'b01010100:  data_out <= 12'b010100101000;
	8'b01010101:  data_out <= 12'b010100101111;
	8'b01010110:  data_out <= 12'b010100110001;
	8'b01010111:  data_out <= 12'b010100110110;
	8'b01011000:  data_out <= 12'b010101001001;
	8'b01011001:  data_out <= 12'b010101001110;
	8'b01011010:  data_out <= 12'b010101010000;
	8'b01011011:  data_out <= 12'b010101010111;
	8'b01011100:  data_out <= 12'b010101100011;
	8'b01011101:  data_out <= 12'b010101100100;
	8'b01011110:  data_out <= 12'b010101111010;
	8'b01011111:  data_out <= 12'b010101111101;
	8'b01100000:  data_out <= 12'b011000000001;
	8'b01100001:  data_out <= 12'b011000000110;
	8'b01100010:  data_out <= 12'b011000011000;
	8'b01100011:  data_out <= 12'b011000011111;
	8'b01100100:  data_out <= 12'b011000101011;
	8'b01100101:  data_out <= 12'b011000101100;
	8'b01100110:  data_out <= 12'b011000110010;
	8'b01100111:  data_out <= 12'b011000110101;
	8'b01101000:  data_out <= 12'b011001001010;
	8'b01101001:  data_out <= 12'b011001001101;
	8'b01101010:  data_out <= 12'b011001010011;
	8'b01101011:  data_out <= 12'b011001010100;
	8'b01101100:  data_out <= 12'b011001100000;
	8'b01101101:  data_out <= 12'b011001100111;
	8'b01101110:  data_out <= 12'b011001111001;
	8'b01101111:  data_out <= 12'b011001111110;
	8'b01110000:  data_out <= 12'b011110000000;
	8'b01110001:  data_out <= 12'b011110000111;
	8'b01110010:  data_out <= 12'b011110011001;
	8'b01110011:  data_out <= 12'b011110011110;
	8'b01110100:  data_out <= 12'b011110101010;
	8'b01110101:  data_out <= 12'b011110101101;
	8'b01110110:  data_out <= 12'b011110110011;
	8'b01110111:  data_out <= 12'b011110110100;
	8'b01111000:  data_out <= 12'b011111001011;
	8'b01111001:  data_out <= 12'b011111001100;
	8'b01111010:  data_out <= 12'b011111010010;
	8'b01111011:  data_out <= 12'b011111010101;
	8'b01111100:  data_out <= 12'b011111100001;
	8'b01111101:  data_out <= 12'b011111100110;
	8'b01111110:  data_out <= 12'b011111111000;
	8'b01111111:  data_out <= 12'b011111111111;
	8'b10000000:  data_out <= 12'b100010001000;
	8'b10000001:  data_out <= 12'b100010001111;
	8'b10000010:  data_out <= 12'b100010010001;
	8'b10000011:  data_out <= 12'b100010010110;
	8'b10000100:  data_out <= 12'b100010100010;
	8'b10000101:  data_out <= 12'b100010100101;
	8'b10000110:  data_out <= 12'b100010111011;
	8'b10000111:  data_out <= 12'b100010111100;
	8'b10001000:  data_out <= 12'b100011000011;
	8'b10001001:  data_out <= 12'b100011000100;
	8'b10001010:  data_out <= 12'b100011011010;
	8'b10001011:  data_out <= 12'b100011011101;
	8'b10001100:  data_out <= 12'b100011101001;
	8'b10001101:  data_out <= 12'b100011101110;
	8'b10001110:  data_out <= 12'b100011110000;
	8'b10001111:  data_out <= 12'b100011110111;
	8'b10010000:  data_out <= 12'b100100001001;
	8'b10010001:  data_out <= 12'b100100001110;
	8'b10010010:  data_out <= 12'b100100010000;
	8'b10010011:  data_out <= 12'b100100010111;
	8'b10010100:  data_out <= 12'b100100100011;
	8'b10010101:  data_out <= 12'b100100100100;
	8'b10010110:  data_out <= 12'b100100111010;
	8'b10010111:  data_out <= 12'b100100111101;
	8'b10011000:  data_out <= 12'b100101000010;
	8'b10011001:  data_out <= 12'b100101000101;
	8'b10011010:  data_out <= 12'b100101011011;
	8'b10011011:  data_out <= 12'b100101011100;
	8'b10011100:  data_out <= 12'b100101101000;
	8'b10011101:  data_out <= 12'b100101101111;
	8'b10011110:  data_out <= 12'b100101110001;
	8'b10011111:  data_out <= 12'b100101110110;
	8'b10100000:  data_out <= 12'b101000001010;
	8'b10100001:  data_out <= 12'b101000001101;
	8'b10100010:  data_out <= 12'b101000010011;
	8'b10100011:  data_out <= 12'b101000010100;
	8'b10100100:  data_out <= 12'b101000100000;
	8'b10100101:  data_out <= 12'b101000100111;
	8'b10100110:  data_out <= 12'b101000111001;
	8'b10100111:  data_out <= 12'b101000111110;
	8'b10101000:  data_out <= 12'b101001000001;
	8'b10101001:  data_out <= 12'b101001000110;
	8'b10101010:  data_out <= 12'b101001011000;
	8'b10101011:  data_out <= 12'b101001011111;
	8'b10101100:  data_out <= 12'b101001101011;
	8'b10101101:  data_out <= 12'b101001101100;
	8'b10101110:  data_out <= 12'b101001110010;
	8'b10101111:  data_out <= 12'b101001110101;
	8'b10110000:  data_out <= 12'b101110001011;
	8'b10110001:  data_out <= 12'b101110001100;
	8'b10110010:  data_out <= 12'b101110010010;
	8'b10110011:  data_out <= 12'b101110010101;
	8'b10110100:  data_out <= 12'b101110100001;
	8'b10110101:  data_out <= 12'b101110100110;
	8'b10110110:  data_out <= 12'b101110111000;
	8'b10110111:  data_out <= 12'b101110111111;
	8'b10111000:  data_out <= 12'b101111000000;
	8'b10111001:  data_out <= 12'b101111000111;
	8'b10111010:  data_out <= 12'b101111011001;
	8'b10111011:  data_out <= 12'b101111011110;
	8'b10111100:  data_out <= 12'b101111101010;
	8'b10111101:  data_out <= 12'b101111101101;
	8'b10111110:  data_out <= 12'b101111110011;
	8'b10111111:  data_out <= 12'b101111110100;
	8'b11000000:  data_out <= 12'b110000001011;
	8'b11000001:  data_out <= 12'b110000001100;
	8'b11000010:  data_out <= 12'b110000010010;
	8'b11000011:  data_out <= 12'b110000010101;
	8'b11000100:  data_out <= 12'b110000100001;
	8'b11000101:  data_out <= 12'b110000100110;
	8'b11000110:  data_out <= 12'b110000111000;
	8'b11000111:  data_out <= 12'b110000111111;
	8'b11001000:  data_out <= 12'b110001000000;
	8'b11001001:  data_out <= 12'b110001000111;
	8'b11001010:  data_out <= 12'b110001011001;
	8'b11001011:  data_out <= 12'b110001011110;
	8'b11001100:  data_out <= 12'b110001101010;
	8'b11001101:  data_out <= 12'b110001101101;
	8'b11001110:  data_out <= 12'b110001110011;
	8'b11001111:  data_out <= 12'b110001110100;
	8'b11010000:  data_out <= 12'b110110001010;
	8'b11010001:  data_out <= 12'b110110001101;
	8'b11010010:  data_out <= 12'b110110010011;
	8'b11010011:  data_out <= 12'b110110010100;
	8'b11010100:  data_out <= 12'b110110100000;
	8'b11010101:  data_out <= 12'b110110100111;
	8'b11010110:  data_out <= 12'b110110111001;
	8'b11010111:  data_out <= 12'b110110111110;
	8'b11011000:  data_out <= 12'b110111000001;
	8'b11011001:  data_out <= 12'b110111000110;
	8'b11011010:  data_out <= 12'b110111011000;
	8'b11011011:  data_out <= 12'b110111011111;
	8'b11011100:  data_out <= 12'b110111101011;
	8'b11011101:  data_out <= 12'b110111101100;
	8'b11011110:  data_out <= 12'b110111110010;
	8'b11011111:  data_out <= 12'b110111110101;
	8'b11100000:  data_out <= 12'b111010001001;
	8'b11100001:  data_out <= 12'b111010001110;
	8'b11100010:  data_out <= 12'b111010010000;
	8'b11100011:  data_out <= 12'b111010010111;
	8'b11100100:  data_out <= 12'b111010100011;
	8'b11100101:  data_out <= 12'b111010100100;
	8'b11100110:  data_out <= 12'b111010111010;
	8'b11100111:  data_out <= 12'b111010111101;
	8'b11101000:  data_out <= 12'b111011000010;
	8'b11101001:  data_out <= 12'b111011000101;
	8'b11101010:  data_out <= 12'b111011011011;
	8'b11101011:  data_out <= 12'b111011011100;
	8'b11101100:  data_out <= 12'b111011101000;
	8'b11101101:  data_out <= 12'b111011101111;
	8'b11101110:  data_out <= 12'b111011110001;
	8'b11101111:  data_out <= 12'b111011110110;
	8'b11110000:  data_out <= 12'b111100001000;
	8'b11110001:  data_out <= 12'b111100001111;
	8'b11110010:  data_out <= 12'b111100010001;
	8'b11110011:  data_out <= 12'b111100010110;
	8'b11110100:  data_out <= 12'b111100100010;
	8'b11110101:  data_out <= 12'b111100100101;
	8'b11110110:  data_out <= 12'b111100111011;
	8'b11110111:  data_out <= 12'b111100111100;
	8'b11111000:  data_out <= 12'b111101000011;
	8'b11111001:  data_out <= 12'b111101000100;
	8'b11111010:  data_out <= 12'b111101011010;
	8'b11111011:  data_out <= 12'b111101011101;
	8'b11111100:  data_out <= 12'b111101101001;
	8'b11111101:  data_out <= 12'b111101101110;
	8'b11111110:  data_out <= 12'b111101110000;
	8'b11111111:  data_out <= 12'b111101110111;
endcase
endmodule
